library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PidController is
  port (
    Clk               : in  std_logic;
    Rst               : in  std_logic
  );
end PidController;

architecture Behavioral of PidController is

begin

end Behavioral;